[info] welcome to sbt 1.10.5 (Eclipse Adoptium Java 17.0.13)
[info] loading project definition from /Users/zach/src/_-genesys2-vivado/keyboard/project
[info] loading settings for project hello from build.sbt ...
[info] set current project to Chisel Example (in build file:/Users/zach/src/_-genesys2-vivado/keyboard/)
[info] compiling 1 Scala source to /Users/zach/src/_-genesys2-vivado/keyboard/target/scala-2.13/classes ...
[info] done compiling
[info] running Main 
// Generated by CIRCT firtool-1.62.1-1-gdf5ed6ea5
// external module IBUFDS

// external module PS2Receiver

// external module Uart_buf_con

// external module Uart_tx

module Top(
  input  clock,
         reset,
         io_PS2Clk,
         io_PS2Data,
  output io_tx
);

  wire        _uart_tx_ready;
  wire        _uart_buf_con_tstart;
  wire [7:0]  _uart_buf_con_tbus;
  wire [15:0] _uut_keycode;
  wire        _uut_oflag;
  reg         start;
  reg  [15:0] keycodev;
  reg  [2:0]  bcount;
  reg         cn;
  reg  [7:0]  keycode_b;
  always @(posedge clock) begin
    if (reset) begin
      start <= 1'h0;
      keycodev <= 16'h0;
      bcount <= 3'h0;
      cn <= 1'h0;
      keycode_b <= 8'h0;
    end
    else begin
      automatic logic _GEN = _uut_oflag & cn;
      start <= _GEN;
      if (_GEN)
        keycodev <= _uut_keycode;
      if (~({8'h0, keycode_b} == _uut_keycode)) begin
        automatic logic _GEN_0 = _uut_keycode[7:0] == 8'hF0;
        automatic logic _GEN_1 = _uut_keycode[15:8] == 8'hF0;
        bcount <= _GEN_0 ? 3'h0 : _GEN_1 ? 3'h5 : 3'h3;
        cn <=
          ~_GEN_0
          & (_GEN_1
               ? _uut_keycode != keycodev
               : {8'h0, _uut_keycode[7:0]} != keycodev | keycodev[15:8] == 8'hF0);
        keycode_b <= _uut_keycode[7:0];
      end
    end
  end // always @(posedge)
  PS2Receiver uut (
    .clk     (clock),
    .kclk    (io_PS2Clk),
    .kdata   (io_PS2Data),
    .keycode (_uut_keycode),
    .oflag   (_uut_oflag)
  );
  Uart_buf_con uart_buf_con (
    .clk    (clock),
    .bcount (bcount),
    .tbuf   (32'h0),
    .start  (start),
    .ready  (/* unused */),
    .tstart (_uart_buf_con_tstart),
    .tready (_uart_tx_ready),
    .tbus   (_uart_buf_con_tbus)
  );
  Uart_tx uart_tx (
    .clk   (clock),
    .tbus  (_uart_buf_con_tbus),
    .start (_uart_buf_con_tstart),
    .tx    (io_tx),
    .ready (_uart_tx_ready)
  );
endmodule

module TopWrapper(
  input  clk_p,
         clk_n,
         reset,
         PS2Data,
         PS2Clk,
  output tx
);

  wire _ibufds_O;
  IBUFDS #(
    .DIFF_TERM("FALSE"),
    .IOSTANDARD("DEFAULT")
  ) ibufds (
    .O  (_ibufds_O),
    .I  (clk_p),
    .IB (clk_n)
  );
  Top top (
    .clock      (_ibufds_O),
    .reset      (reset),
    .io_PS2Clk  (PS2Clk),
    .io_PS2Data (PS2Data),
    .io_tx      (tx)
  );
endmodule


// ----- 8< ----- FILE "./PS2Receiver.v" ----- 8< -----

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Digilent Inc.
// Engineer: Thomas Kappenman
//
// Create Date: 03/03/2015 09:33:36 PM
// Design Name:
// Module Name: PS2Receiver
// Project Name: Nexys4DDR Keyboard Demo
// Target Devices: Nexys4DDR
// Tool Versions:
// Description: PS2 Receiver module used to shift in keycodes from a keyboard plugged into the PS2 port
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module PS2Receiver(
    input clk,
    input kclk,
    input kdata,
    output reg [15:0] keycode=0,
    output reg oflag
    );

    wire kclkf, kdataf;
    reg [7:0]datacur=0;
    reg [7:0]dataprev=0;
    reg [3:0]cnt=0;
    reg flag=0;

debouncer #(
    .COUNT_MAX(76),
    .COUNT_WIDTH(7)
) db_clk(
    .clk(clk),
    .I(kclk),
    .O(kclkf)
);
debouncer #(
   .COUNT_MAX(76),
   .COUNT_WIDTH(7)
) db_data(
    .clk(clk),
    .I(kdata),
    .O(kdataf)
);

always@(negedge(kclkf))begin
    case(cnt)
    0:;//Start bit
    1:datacur[0]<=kdataf;
    2:datacur[1]<=kdataf;
    3:datacur[2]<=kdataf;
    4:datacur[3]<=kdataf;
    5:datacur[4]<=kdataf;
    6:datacur[5]<=kdataf;
    7:datacur[6]<=kdataf;
    8:datacur[7]<=kdataf;
    9:flag<=1'b1;
    10:flag<=1'b0;

    endcase
        if(cnt<=9) cnt<=cnt+1;
        else if(cnt==10) cnt<=0;
end

reg pflag;
always@(posedge clk) begin
    if (flag == 1'b1 && pflag == 1'b0) begin
        keycode <= {dataprev, datacur};
        oflag <= 1'b1;
        dataprev <= datacur;
    end else
        oflag <= 'b0;
    pflag <= flag;
end

endmodule

// ----- 8< ----- FILE "./debouncer.v" ----- 8< -----

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 07/27/2016 02:04:22 PM
// Design Name:
// Module Name: debouncer
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module debouncer(
    input clk,
    input I,
    output reg O
    );
    parameter COUNT_MAX=255, COUNT_WIDTH=8;
    reg [COUNT_WIDTH-1:0] count;
    reg Iv=0;
    always@(posedge clk)
        if (I == Iv) begin
            if (count == COUNT_MAX)
                O <= I;
            else
                count <= count + 1'b1;
        end else begin
            count <= 'b0;
            Iv <= I;
        end

endmodule

// ----- 8< ----- FILE "./uart_buf_con.v" ----- 8< -----

module uart_buf_con(
    input             clk,
    input      [ 2:0] bcount,
    input      [31:0] tbuf,
    input             start,
    output            ready,
    output reg        tstart=0,
    input             tready,
    output reg [ 7:0] tbus=0
    );
    reg [2:0] sel=0;
    reg [31:0] pbuf=0;
    reg running=0;
    initial tstart <= 'b0;
    initial tbus <= 'b0;
    always@(posedge clk)
        if (tready == 1'b1) begin
            if (running == 1'b1) begin
                if (sel == 4'd1) begin
                    running <= 1'b0;
                    sel <= bcount + 2'd2;
                end else begin
                    sel <= sel - 1'b1;
                    tstart <= 1'b1;
                    running <= 1'b1;
                end
            end else begin
                if (bcount != 2'b0) begin
                    pbuf <= tbuf;
                    tstart <= start;
                    running <= start;
                    sel <= bcount + 2'd2;
                end
            end
        end else
            tstart <= 1'b0;
    assign ready = ~running;
    always@(sel, pbuf)
        case (sel)
        1: tbus <= 8'd13;
        2: tbus <= 8'd10;
        3: tbus <= pbuf[7:0];
        4: tbus <= pbuf[15:8];
        5: tbus <= 8'd32;
        6: tbus <= pbuf[23:16];
        7: tbus <= pbuf[31:24];
        default: tbus <= 8'd0;
        endcase
endmodule

// ----- 8< ----- FILE "./uart_tx.v" ----- 8< -----


module uart_tx(
    input       clk   ,
    input [7:0] tbus  ,
    input       start,
    output      tx    ,
    output      ready
    );
    parameter CD_MAX=10416, CD_WIDTH=16;
    reg [CD_WIDTH-1:0] cd_count=0;
    reg [3:0] count=0;
    reg running=0;
    reg [10:0] shift=11'h7ff;
    always@(posedge clk) begin
        if (running == 1'b0) begin
            shift <= {2'b11, tbus, 1'b0};
            running <= start;
            cd_count <= 'b0;
            count <= 'b0;
        end else if (cd_count == CD_MAX) begin
            shift <= {1'b1, shift[10:1]};
            cd_count <= 'b0;
            if (count == 4'd10) begin
                running <= 1'b0;
                count <= 'b0;
            end
            else
                count <= count + 1'b1;
        end else
            cd_count <= cd_count + 1'b1;
    end
    assign tx = (running == 1'b1) ? shift[0] : 1'b1;
    assign ready = ((running == 1'b0 && start == 1'b0) || (cd_count == CD_MAX && count == 4'd10)) ? 1'b1 : 1'b0;
endmodule

// ----- 8< ----- FILE "firrtl_black_box_resource_files.f" ----- 8< -----

PS2Receiver.v
debouncer.v
uart_buf_con.v
uart_tx.v

[success] Total time: 4 s, completed Dec 10, 2024, 1:09:15 PM
